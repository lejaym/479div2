magic
tech scmos
timestamp 1428619208
<< pwell >>
rect 993 1561 1103 1570
rect 993 1548 1653 1561
rect 993 1542 1213 1548
rect 1103 1515 1213 1542
rect 1103 1370 1213 1426
rect 1425 1370 1438 1380
rect 902 1185 926 1267
rect 1103 1169 1213 1251
rect 1727 986 1773 1068
<< nwell >>
rect 1103 1432 1213 1509
rect 1103 1257 1213 1364
rect 903 1121 926 1181
rect 909 1116 926 1121
rect 1103 1115 1213 1163
rect 1711 1071 1773 1117
<< polysilicon >>
rect 1125 1525 1127 1527
rect 1137 1525 1163 1527
rect 1159 1523 1163 1525
rect 1177 1525 1180 1527
rect 1190 1525 1204 1527
rect 1159 1500 1167 1523
rect 1125 1498 1127 1500
rect 1147 1498 1156 1500
rect 1159 1498 1170 1500
rect 1190 1498 1192 1500
rect 1151 1489 1156 1498
rect 1151 1483 1161 1489
rect 1125 1459 1127 1461
rect 1177 1459 1179 1461
rect 1125 1437 1127 1439
rect 1177 1437 1179 1439
rect 1114 1435 1127 1437
rect 1121 1425 1127 1435
rect 1114 1423 1127 1425
rect 1157 1435 1179 1437
rect 1164 1425 1179 1435
rect 1707 1433 1715 1434
rect 1157 1423 1179 1425
rect 1125 1421 1127 1423
rect 1177 1421 1179 1423
rect 1125 1409 1127 1411
rect 1177 1409 1179 1411
rect 1148 1386 1150 1388
rect 1185 1386 1187 1388
rect 1148 1374 1150 1376
rect 1148 1372 1165 1374
rect 1148 1362 1158 1372
rect 1148 1360 1165 1362
rect 1185 1372 1187 1376
rect 1185 1370 1210 1372
rect 1185 1364 1197 1370
rect 1185 1362 1210 1364
rect 1148 1358 1150 1360
rect 1185 1358 1187 1362
rect 1148 1336 1150 1338
rect 1185 1336 1187 1338
rect 1710 1329 1712 1433
rect 1730 1410 1732 1434
rect 1740 1410 1742 1434
rect 1730 1328 1732 1365
rect 1740 1329 1742 1362
rect 1168 1312 1170 1314
rect 1193 1312 1195 1314
rect 1118 1276 1125 1311
rect 1128 1292 1130 1294
rect 1150 1292 1159 1294
rect 1118 1274 1130 1276
rect 1150 1274 1152 1276
rect 1118 1235 1125 1274
rect 1154 1253 1159 1292
rect 1168 1271 1170 1273
rect 1179 1271 1184 1297
rect 1193 1290 1195 1292
rect 1193 1287 1208 1290
rect 1193 1283 1195 1285
rect 1168 1264 1184 1271
rect 1153 1245 1159 1253
rect 1128 1243 1130 1245
rect 1140 1243 1159 1245
rect 1179 1259 1184 1264
rect 1193 1259 1195 1263
rect 1179 1249 1195 1259
rect 1118 1233 1128 1235
rect 1126 1227 1128 1233
rect 1126 1225 1130 1227
rect 1140 1225 1143 1227
rect 1179 1226 1184 1249
rect 1193 1247 1195 1249
rect 1193 1235 1195 1237
rect 1203 1233 1208 1287
rect 1193 1229 1208 1233
rect 1193 1227 1195 1229
rect 1203 1226 1208 1229
rect 1193 1215 1195 1217
rect 912 1198 914 1200
rect 912 1178 914 1188
rect 1136 1185 1138 1187
rect 1178 1185 1180 1187
rect 1136 1173 1138 1175
rect 1178 1173 1180 1175
rect 1136 1171 1153 1173
rect 1136 1161 1146 1171
rect 1136 1159 1153 1161
rect 1178 1171 1191 1173
rect 1178 1161 1184 1171
rect 1178 1159 1191 1161
rect 912 1156 914 1158
rect 1136 1157 1138 1159
rect 1178 1157 1180 1159
rect 1136 1135 1138 1137
rect 1178 1135 1180 1137
rect 1754 1097 1755 1101
rect 1735 1093 1737 1095
rect 1753 1093 1755 1097
rect 1763 1097 1764 1101
rect 1763 1093 1765 1097
rect 1735 1072 1737 1075
rect 1735 1068 1736 1072
rect 1735 1065 1737 1068
rect 1753 1065 1755 1075
rect 1763 1065 1765 1075
rect 1735 1053 1737 1055
rect 1753 1053 1755 1055
rect 1763 1053 1765 1055
<< ndiffusion >>
rect 1127 1527 1137 1528
rect 1127 1524 1137 1525
rect 1180 1527 1190 1528
rect 1180 1524 1190 1525
rect 1124 1411 1125 1421
rect 1127 1411 1128 1421
rect 1176 1411 1177 1421
rect 1179 1411 1180 1421
rect 1147 1376 1148 1386
rect 1150 1376 1151 1386
rect 1184 1376 1185 1386
rect 1187 1376 1188 1386
rect 1130 1245 1140 1246
rect 1130 1242 1140 1243
rect 1130 1227 1140 1228
rect 1192 1237 1193 1247
rect 1195 1237 1196 1247
rect 1130 1224 1140 1225
rect 1192 1217 1193 1227
rect 1195 1217 1196 1227
rect 910 1188 912 1198
rect 914 1188 916 1198
rect 1135 1175 1136 1185
rect 1138 1175 1139 1185
rect 1177 1175 1178 1185
rect 1180 1175 1181 1185
rect 1733 1055 1735 1065
rect 1737 1055 1739 1065
rect 1751 1055 1753 1065
rect 1755 1055 1757 1065
rect 1761 1055 1763 1065
rect 1765 1055 1767 1065
<< pdiffusion >>
rect 1127 1500 1147 1501
rect 1170 1500 1190 1501
rect 1127 1497 1147 1498
rect 1170 1497 1190 1498
rect 1124 1439 1125 1459
rect 1127 1439 1128 1459
rect 1176 1439 1177 1459
rect 1179 1439 1180 1459
rect 1147 1338 1148 1358
rect 1150 1338 1151 1358
rect 1184 1338 1185 1358
rect 1187 1338 1188 1358
rect 1130 1294 1150 1295
rect 1130 1291 1150 1292
rect 1130 1276 1150 1277
rect 1130 1273 1150 1274
rect 1167 1273 1168 1312
rect 1170 1273 1171 1312
rect 1192 1292 1193 1312
rect 1195 1292 1196 1312
rect 1192 1263 1193 1283
rect 1195 1263 1196 1283
rect 910 1158 912 1178
rect 914 1158 916 1178
rect 1135 1137 1136 1157
rect 1138 1137 1139 1157
rect 1177 1137 1178 1157
rect 1180 1137 1181 1157
rect 1733 1075 1735 1093
rect 1737 1075 1739 1093
rect 1751 1075 1753 1093
rect 1755 1075 1757 1093
rect 1761 1075 1763 1093
rect 1765 1075 1767 1093
<< metal1 >>
rect 870 2018 1715 2026
rect 870 1888 878 2018
rect 928 2006 1704 2014
rect 20 1880 878 1888
rect 882 1984 998 2000
rect 1645 1984 1689 2000
rect 882 1876 916 1984
rect 1420 1946 1434 1952
rect -36 1840 916 1876
rect 938 1910 1001 1926
rect -35 1778 5 1840
rect 43 1821 49 1828
rect 938 1823 976 1910
rect 910 1807 976 1823
rect -34 1749 4 1778
rect -34 1733 30 1749
rect -34 1560 4 1733
rect 938 1725 976 1807
rect 1665 1799 1689 1984
rect 1642 1783 1689 1799
rect 1424 1742 1430 1751
rect 938 1709 1001 1725
rect 938 1675 976 1709
rect 909 1659 976 1675
rect 915 1635 920 1643
rect 910 1617 917 1623
rect 938 1577 976 1659
rect 1665 1651 1689 1783
rect 1642 1635 1689 1651
rect 938 1561 1000 1577
rect -34 1544 30 1560
rect 938 1554 1653 1561
rect -34 1359 4 1544
rect 938 1538 1002 1554
rect 1103 1552 1213 1554
rect 1103 1540 1117 1552
rect 1124 1540 1145 1552
rect 1152 1540 1174 1552
rect 1181 1540 1213 1552
rect 1103 1538 1213 1540
rect 910 1446 929 1454
rect 938 1433 976 1538
rect 1116 1528 1127 1532
rect 1116 1516 1124 1528
rect 1116 1510 1118 1516
rect 1116 1497 1124 1510
rect 1152 1523 1163 1529
rect 1190 1528 1200 1532
rect 1127 1516 1190 1520
rect 1127 1510 1131 1516
rect 1137 1510 1190 1516
rect 1127 1505 1190 1510
rect 1193 1515 1200 1528
rect 1199 1509 1200 1515
rect 1193 1497 1200 1509
rect 1116 1493 1127 1497
rect 1190 1493 1200 1497
rect 1167 1484 1172 1489
rect 1204 1489 1210 1523
rect 1178 1484 1210 1489
rect 1167 1483 1210 1484
rect 1103 1478 1213 1480
rect 1103 1466 1119 1478
rect 1126 1466 1144 1478
rect 1151 1466 1182 1478
rect 1189 1466 1213 1478
rect 1336 1477 1344 1494
rect 1665 1480 1689 1635
rect 1103 1464 1213 1466
rect 1642 1464 1647 1480
rect 1654 1464 1689 1480
rect 1116 1459 1124 1464
rect 1168 1459 1176 1464
rect 1116 1439 1120 1459
rect 1132 1439 1152 1459
rect 1168 1439 1172 1459
rect 1184 1439 1201 1459
rect 1140 1437 1152 1439
rect 1140 1435 1164 1437
rect 910 1417 976 1433
rect 1121 1433 1136 1435
rect 1121 1427 1130 1433
rect 1121 1425 1136 1427
rect 1140 1425 1157 1435
rect 1140 1423 1164 1425
rect 1189 1434 1201 1439
rect 1189 1428 1190 1434
rect 1196 1428 1201 1434
rect 1140 1421 1152 1423
rect 1189 1421 1201 1428
rect 938 1406 976 1417
rect 1116 1411 1120 1421
rect 1132 1420 1152 1421
rect 1132 1413 1136 1420
rect 1143 1413 1152 1420
rect 1132 1411 1152 1413
rect 1168 1411 1172 1421
rect 1184 1411 1201 1421
rect 1675 1418 1689 1464
rect 1696 1431 1704 2006
rect 1707 1442 1715 2018
rect 1696 1423 1764 1431
rect 1675 1414 1711 1418
rect 1116 1406 1124 1411
rect 1168 1406 1176 1411
rect 938 1390 999 1406
rect 1103 1404 1213 1406
rect 1103 1392 1117 1404
rect 1124 1392 1145 1404
rect 1152 1392 1174 1404
rect 1181 1392 1213 1404
rect 1103 1390 1213 1392
rect 1655 1390 1670 1406
rect 1682 1398 1707 1411
rect -34 1339 30 1359
rect -34 1124 4 1339
rect 938 1229 976 1390
rect 1151 1386 1159 1390
rect 1188 1386 1196 1390
rect 1138 1372 1143 1386
rect 1155 1376 1159 1386
rect 1165 1376 1180 1386
rect 1192 1376 1196 1386
rect 1661 1381 1688 1390
rect 1699 1387 1707 1398
rect 1699 1383 1711 1387
rect 1103 1362 1143 1372
rect 1128 1361 1143 1362
rect 1128 1355 1135 1361
rect 1141 1355 1143 1361
rect 1165 1358 1177 1376
rect 1424 1372 1433 1375
rect 1203 1370 1213 1372
rect 1427 1371 1433 1372
rect 1210 1364 1213 1370
rect 1203 1362 1213 1364
rect 1671 1363 1680 1372
rect 1684 1366 1688 1381
rect 1684 1362 1712 1366
rect 1128 1338 1143 1355
rect 1155 1338 1159 1358
rect 1165 1349 1180 1358
rect 1165 1342 1169 1349
rect 1176 1342 1180 1349
rect 1165 1338 1180 1342
rect 1192 1338 1196 1358
rect 1756 1348 1764 1423
rect 1151 1332 1159 1338
rect 1188 1332 1196 1338
rect 1103 1330 1213 1332
rect 1103 1319 1119 1330
rect 1126 1319 1144 1330
rect 1151 1319 1182 1330
rect 1189 1319 1213 1330
rect 1103 1316 1213 1319
rect 1171 1312 1175 1316
rect 1196 1312 1200 1316
rect 1779 1314 1824 1318
rect 1133 1305 1137 1311
rect 1113 1295 1130 1299
rect 1113 1239 1119 1295
rect 1150 1287 1163 1291
rect 1130 1281 1163 1287
rect 1150 1277 1163 1281
rect 1125 1269 1130 1273
rect 1125 1262 1140 1269
rect 1125 1255 1131 1262
rect 1138 1255 1140 1262
rect 1125 1250 1140 1255
rect 1125 1246 1130 1250
rect 1151 1259 1153 1265
rect 1145 1253 1153 1259
rect 1145 1245 1148 1253
rect 1156 1260 1163 1277
rect 1179 1308 1188 1312
rect 1184 1297 1188 1308
rect 1179 1292 1188 1297
rect 1196 1283 1200 1292
rect 1775 1291 1793 1295
rect 1156 1253 1175 1260
rect 1156 1247 1169 1253
rect 1113 1234 1125 1239
rect 910 1221 976 1229
rect 1117 1226 1125 1234
rect 1156 1238 1163 1247
rect 1183 1241 1188 1283
rect 1779 1260 1786 1264
rect 1130 1232 1163 1238
rect 1167 1232 1188 1241
rect 916 1198 920 1221
rect 938 1205 976 1221
rect 991 1218 999 1226
rect 1103 1218 1114 1226
rect 1123 1224 1125 1226
rect 1123 1220 1130 1224
rect 1108 1216 1114 1218
rect 1167 1216 1175 1232
rect 1196 1227 1200 1237
rect 1179 1226 1188 1227
rect 1184 1218 1188 1226
rect 1179 1217 1188 1218
rect 1209 1218 1213 1226
rect 1108 1208 1175 1216
rect 1196 1205 1200 1217
rect 938 1189 998 1205
rect 1103 1203 1213 1205
rect 1103 1191 1117 1203
rect 1124 1191 1145 1203
rect 1152 1191 1174 1203
rect 1181 1191 1213 1203
rect 1103 1189 1213 1191
rect 1778 1189 1786 1193
rect 906 1178 910 1188
rect 918 1181 921 1185
rect 916 1124 920 1158
rect -34 1116 30 1124
rect 907 1116 920 1124
rect -34 893 4 1116
rect 20 1022 48 1039
rect 938 1021 976 1189
rect 1139 1185 1147 1189
rect 1181 1185 1189 1189
rect 1114 1175 1131 1185
rect 1143 1175 1147 1185
rect 1153 1175 1173 1185
rect 1185 1175 1189 1185
rect 1114 1168 1126 1175
rect 1114 1162 1119 1168
rect 1125 1162 1126 1168
rect 1114 1157 1126 1162
rect 1153 1157 1165 1175
rect 1169 1169 1184 1171
rect 1175 1163 1184 1169
rect 1169 1161 1184 1163
rect 1114 1137 1131 1157
rect 1143 1137 1147 1157
rect 1153 1148 1173 1157
rect 1153 1141 1157 1148
rect 1164 1141 1173 1148
rect 1153 1137 1173 1141
rect 1185 1137 1189 1157
rect 1139 1131 1147 1137
rect 1181 1131 1189 1137
rect 1103 1129 1213 1131
rect 1103 1117 1119 1129
rect 1126 1117 1144 1129
rect 1151 1117 1182 1129
rect 1189 1117 1213 1129
rect 1103 1115 1213 1117
rect 1743 1115 1746 1116
rect 1743 1100 1747 1115
rect 1739 1096 1747 1100
rect 1750 1101 1754 1105
rect 1739 1093 1743 1096
rect 1757 1093 1761 1117
rect 1768 1097 1772 1101
rect 1729 1065 1733 1075
rect 1747 1072 1751 1075
rect 1767 1072 1771 1075
rect 1740 1068 1771 1072
rect 1747 1065 1751 1068
rect 987 1049 1513 1052
rect 1729 1049 1733 1055
rect 987 1044 1733 1049
rect 1739 1044 1743 1055
rect 1767 1044 1771 1055
rect 1739 1040 1771 1044
rect 987 1028 1744 1036
rect 1755 1021 1759 1040
rect 1782 1036 1786 1189
rect 1789 1101 1793 1291
rect 1770 1028 1786 1036
rect 1796 1028 1800 1256
rect 1804 1028 1808 1264
rect 1812 1028 1816 1158
rect 1820 1028 1824 1314
rect 1828 1028 1836 1105
rect 1844 1028 1852 1048
rect 938 998 1865 1021
rect 910 997 1865 998
rect 909 993 1865 997
rect 1785 986 1865 993
rect -34 878 30 893
rect -34 670 4 878
rect 1828 785 1865 986
rect 1787 769 1865 785
rect 1795 745 1796 753
rect 1790 727 1804 733
rect -34 654 30 670
rect -34 524 4 654
rect 1828 555 1865 769
rect 1790 547 1865 555
rect -34 513 30 524
rect -34 385 4 513
rect 1828 459 1865 547
rect 1787 443 1865 459
rect -34 369 30 385
rect -34 237 4 369
rect 1828 311 1865 443
rect 1790 295 1865 311
rect 1790 267 1798 277
rect -34 220 30 237
rect -34 36 4 220
rect 1790 123 1798 131
rect 1828 110 1865 295
rect 1790 94 1865 110
rect -34 20 31 36
rect 1828 19 1865 94
<< metal2 >>
rect 12 1039 20 1880
rect 43 1833 49 1864
rect 43 1823 49 1828
rect 153 1834 159 1864
rect 153 1823 159 1829
rect 263 1833 269 1864
rect 263 1823 269 1828
rect 373 1834 379 1864
rect 373 1823 379 1829
rect 483 1834 489 1864
rect 483 1823 489 1829
rect 593 1833 599 1864
rect 593 1823 599 1828
rect 703 1833 709 1864
rect 703 1823 709 1828
rect 813 1833 819 1864
rect 813 1823 819 1828
rect 920 1643 928 2006
rect 1056 1984 1110 1990
rect 1163 1984 1220 1990
rect 1275 1984 1330 1990
rect 1387 1984 1420 1990
rect 1496 1984 1550 1990
rect 1594 1986 1607 2029
rect 976 1643 989 1753
rect 925 1635 928 1643
rect 917 1336 925 1617
rect 1104 1605 1110 1984
rect 1214 1605 1220 1984
rect 1324 1605 1330 1984
rect 1414 1952 1420 1984
rect 1104 1599 1124 1605
rect 1214 1599 1229 1605
rect 1324 1599 1344 1605
rect 995 1565 1011 1571
rect 935 1446 991 1454
rect 917 1328 949 1336
rect 910 1316 933 1320
rect 925 1036 933 1316
rect 941 1052 949 1328
rect 981 1226 991 1446
rect 995 1132 1001 1565
rect 1118 1550 1124 1552
rect 1010 1544 1113 1550
rect 1107 1132 1113 1544
rect 1118 1544 1223 1550
rect 1118 1516 1124 1544
rect 1149 1535 1159 1536
rect 1149 1529 1152 1535
rect 1158 1529 1159 1535
rect 1128 1516 1139 1517
rect 1128 1510 1131 1516
rect 1137 1510 1139 1516
rect 1128 1433 1139 1510
rect 1128 1427 1130 1433
rect 1136 1427 1139 1433
rect 1128 1426 1139 1427
rect 1121 1420 1143 1422
rect 1121 1413 1136 1420
rect 1121 1411 1143 1413
rect 1121 1264 1128 1411
rect 1149 1397 1159 1529
rect 1188 1509 1193 1515
rect 1135 1390 1159 1397
rect 1167 1484 1172 1490
rect 1135 1361 1144 1390
rect 1141 1355 1144 1361
rect 1135 1311 1144 1355
rect 1167 1349 1178 1484
rect 1188 1434 1199 1509
rect 1188 1428 1190 1434
rect 1196 1428 1199 1434
rect 1188 1426 1199 1428
rect 1167 1342 1169 1349
rect 1176 1342 1178 1349
rect 1167 1341 1178 1342
rect 1135 1305 1137 1311
rect 1143 1305 1144 1311
rect 1135 1303 1144 1305
rect 1158 1332 1178 1341
rect 1158 1267 1168 1332
rect 1144 1265 1168 1267
rect 1121 1262 1140 1264
rect 1121 1255 1131 1262
rect 1138 1255 1140 1262
rect 1144 1259 1145 1265
rect 1151 1259 1168 1265
rect 1144 1258 1168 1259
rect 1121 1253 1140 1255
rect 1167 1247 1169 1253
rect 1175 1247 1177 1253
rect 1123 1220 1128 1226
rect 1119 1168 1128 1220
rect 1125 1162 1128 1168
rect 1167 1169 1177 1247
rect 1167 1163 1169 1169
rect 1175 1163 1177 1169
rect 1167 1162 1177 1163
rect 1154 1148 1167 1151
rect 1154 1141 1157 1148
rect 1164 1141 1167 1148
rect 1154 1132 1167 1141
rect 995 1126 1055 1132
rect 1107 1126 1167 1132
rect 1217 1132 1223 1544
rect 1229 1542 1333 1548
rect 1327 1133 1333 1542
rect 1424 1381 1430 1731
rect 1434 1605 1440 1946
rect 1544 1605 1550 1984
rect 1661 1889 1696 1897
rect 1661 1743 1682 1753
rect 1434 1599 1454 1605
rect 1544 1599 1564 1605
rect 1647 1332 1654 1464
rect 1674 1411 1682 1743
rect 1686 1348 1696 1889
rect 1653 1316 1673 1332
rect 1786 1264 1804 1268
rect 1778 1256 1796 1260
rect 1778 1158 1812 1162
rect 1755 1135 1865 1139
rect 1217 1126 1268 1132
rect 1327 1127 1385 1133
rect 1154 1115 1167 1126
rect 1754 1105 1828 1112
rect 1779 1097 1789 1101
rect 1005 1088 1869 1092
rect 941 1044 979 1052
rect 925 1028 979 1036
rect 1005 994 1011 1088
rect 1115 1080 1869 1084
rect 1115 994 1121 1080
rect 1225 1072 1869 1076
rect 1225 994 1231 1072
rect 1335 1064 1869 1068
rect 1335 994 1341 1064
rect 1445 1056 1869 1060
rect 1445 994 1451 1056
rect 1555 1048 1869 1052
rect 1555 994 1561 1048
rect 1665 1040 1869 1044
rect 1665 994 1671 1040
rect 1752 1028 1762 1036
rect 1774 1032 1869 1036
rect 1774 994 1780 1032
rect 1796 753 1800 1024
rect 1804 733 1808 1024
rect 1812 501 1816 1024
rect 1790 493 1812 501
rect 1820 469 1824 1024
rect 1790 466 1820 469
rect 1794 462 1820 466
rect 1828 277 1836 1024
rect 1806 267 1836 277
rect 1844 131 1852 1024
rect 1804 123 1852 131
rect 81 17 94 20
rect 81 -21 94 11
rect 191 17 204 20
rect 191 -21 204 11
rect 301 17 314 20
rect 301 -21 314 11
rect 411 17 424 20
rect 411 -21 424 11
rect 521 17 534 20
rect 521 -21 534 11
rect 631 17 644 20
rect 631 -21 644 11
rect 741 17 754 20
rect 741 -21 754 11
rect 851 17 864 20
rect 851 -21 864 11
rect 961 17 974 20
rect 961 -21 974 11
rect 1071 17 1084 20
rect 1071 -21 1084 11
rect 1181 17 1194 20
rect 1181 -21 1194 11
rect 1291 17 1304 20
rect 1291 -21 1304 11
rect 1401 17 1414 20
rect 1401 -21 1414 11
rect 1511 17 1524 20
rect 1511 -21 1524 11
rect 1621 17 1634 20
rect 1621 -21 1634 11
rect 1731 17 1744 20
rect 1731 -21 1744 11
<< ntransistor >>
rect 1127 1525 1137 1527
rect 1180 1525 1190 1527
rect 1125 1411 1127 1421
rect 1177 1411 1179 1421
rect 1148 1376 1150 1386
rect 1185 1376 1187 1386
rect 1130 1243 1140 1245
rect 1130 1225 1140 1227
rect 1193 1237 1195 1247
rect 1193 1217 1195 1227
rect 912 1188 914 1198
rect 1136 1175 1138 1185
rect 1178 1175 1180 1185
rect 1735 1055 1737 1065
rect 1753 1055 1755 1065
rect 1763 1055 1765 1065
<< ptransistor >>
rect 1127 1498 1147 1500
rect 1170 1498 1190 1500
rect 1125 1439 1127 1459
rect 1177 1439 1179 1459
rect 1148 1338 1150 1358
rect 1185 1338 1187 1358
rect 1130 1292 1150 1294
rect 1130 1274 1150 1276
rect 1168 1273 1170 1312
rect 1193 1292 1195 1312
rect 1193 1263 1195 1283
rect 912 1158 914 1178
rect 1136 1137 1138 1157
rect 1178 1137 1180 1157
rect 1735 1075 1737 1093
rect 1753 1075 1755 1093
rect 1763 1075 1765 1093
<< polycontact >>
rect 910 1635 915 1643
rect 1163 1523 1169 1529
rect 1204 1523 1210 1529
rect 1161 1483 1167 1489
rect 1114 1425 1121 1435
rect 1157 1425 1164 1435
rect 1707 1434 1715 1442
rect 1158 1362 1165 1372
rect 1197 1364 1210 1370
rect 1125 1305 1133 1311
rect 1179 1297 1184 1308
rect 1148 1245 1153 1253
rect 1179 1218 1184 1226
rect 1203 1218 1209 1226
rect 914 1181 918 1185
rect 1146 1161 1153 1171
rect 1184 1161 1191 1171
rect 1750 1097 1754 1101
rect 1764 1097 1768 1101
rect 1736 1068 1740 1072
rect 1790 745 1795 753
<< ndcontact >>
rect 1127 1528 1137 1532
rect 1127 1520 1137 1524
rect 1180 1528 1190 1532
rect 1180 1520 1190 1524
rect 1120 1411 1124 1421
rect 1128 1411 1132 1421
rect 1172 1411 1176 1421
rect 1180 1411 1184 1421
rect 1143 1376 1147 1386
rect 1151 1376 1155 1386
rect 1180 1376 1184 1386
rect 1188 1376 1192 1386
rect 1130 1246 1140 1250
rect 1130 1238 1140 1242
rect 1130 1228 1140 1232
rect 1188 1237 1192 1247
rect 1196 1237 1200 1247
rect 1130 1220 1140 1224
rect 1188 1217 1192 1227
rect 1196 1217 1200 1227
rect 906 1188 910 1198
rect 916 1188 920 1198
rect 1131 1175 1135 1185
rect 1139 1175 1143 1185
rect 1173 1175 1177 1185
rect 1181 1175 1185 1185
rect 1729 1055 1733 1065
rect 1739 1055 1743 1065
rect 1747 1055 1751 1065
rect 1757 1055 1761 1065
rect 1767 1055 1771 1065
<< pdcontact >>
rect 1127 1501 1147 1505
rect 1170 1501 1190 1505
rect 1127 1493 1147 1497
rect 1170 1493 1190 1497
rect 1120 1439 1124 1459
rect 1128 1439 1132 1459
rect 1172 1439 1176 1459
rect 1180 1439 1184 1459
rect 1143 1338 1147 1358
rect 1151 1338 1155 1358
rect 1180 1338 1184 1358
rect 1188 1338 1192 1358
rect 1130 1295 1150 1299
rect 1130 1287 1150 1291
rect 1130 1277 1150 1281
rect 1130 1269 1150 1273
rect 1163 1273 1167 1312
rect 1171 1273 1175 1312
rect 1188 1292 1192 1312
rect 1196 1292 1200 1312
rect 1188 1263 1192 1283
rect 1196 1263 1200 1283
rect 906 1158 910 1178
rect 916 1158 920 1178
rect 1131 1137 1135 1157
rect 1139 1137 1143 1157
rect 1173 1137 1177 1157
rect 1181 1137 1185 1157
rect 1729 1075 1733 1093
rect 1739 1075 1743 1093
rect 1747 1075 1751 1093
rect 1757 1075 1761 1093
rect 1767 1075 1771 1093
<< m2contact >>
rect 1594 2029 1607 2033
rect 920 2006 928 2014
rect 12 1880 20 1888
rect 1414 1946 1420 1952
rect 1434 1946 1440 1952
rect 43 1828 49 1833
rect 153 1829 159 1834
rect 263 1828 269 1833
rect 373 1829 379 1834
rect 483 1829 489 1834
rect 593 1828 599 1833
rect 703 1828 709 1833
rect 813 1828 819 1833
rect 1651 1889 1661 1897
rect 989 1743 1002 1753
rect 1651 1743 1661 1753
rect 1424 1731 1430 1742
rect 920 1635 925 1643
rect 917 1617 925 1623
rect 929 1446 935 1454
rect 1152 1529 1158 1535
rect 1118 1510 1124 1516
rect 1131 1510 1137 1516
rect 1193 1509 1199 1515
rect 1172 1484 1178 1490
rect 1647 1464 1654 1480
rect 1130 1427 1136 1433
rect 1190 1428 1196 1434
rect 1136 1413 1143 1420
rect 1674 1398 1682 1411
rect 904 1316 910 1320
rect 1135 1355 1141 1361
rect 1424 1375 1430 1381
rect 1169 1342 1176 1349
rect 1844 1344 1852 1352
rect 1640 1316 1653 1332
rect 1137 1305 1143 1311
rect 1131 1255 1138 1262
rect 1145 1259 1151 1265
rect 1169 1247 1175 1253
rect 1782 1264 1786 1268
rect 981 1218 991 1226
rect 1117 1220 1123 1226
rect 921 1181 925 1185
rect 12 1022 20 1039
rect 1119 1162 1125 1168
rect 1169 1163 1175 1169
rect 1157 1141 1164 1148
rect 1751 1135 1755 1139
rect 1750 1105 1754 1112
rect 1772 1097 1779 1101
rect 979 1044 987 1052
rect 979 1028 987 1036
rect 1744 1028 1752 1036
rect 1804 1264 1808 1268
rect 1789 1097 1793 1101
rect 1796 1256 1800 1260
rect 1762 1028 1770 1036
rect 1796 1024 1800 1028
rect 1804 1024 1808 1028
rect 1812 1158 1816 1162
rect 1812 1024 1816 1028
rect 1820 1024 1824 1028
rect 1828 1105 1836 1112
rect 1828 1024 1836 1028
rect 1844 1024 1852 1028
rect 1796 745 1800 753
rect 1804 727 1808 733
rect 1812 493 1816 501
rect 1790 462 1794 466
rect 1820 462 1824 469
rect 1798 267 1806 277
rect 1798 123 1804 131
rect 81 11 94 17
rect 191 11 204 17
rect 301 11 314 17
rect 411 11 424 17
rect 521 11 534 17
rect 631 11 644 17
rect 741 11 754 17
rect 851 11 864 17
rect 961 11 974 17
rect 1071 11 1084 17
rect 1181 11 1194 17
rect 1291 11 1304 17
rect 1401 11 1414 17
rect 1511 11 1524 17
rect 1621 11 1634 17
rect 1731 11 1744 17
<< psubstratepcontact >>
rect 1117 1540 1124 1552
rect 1145 1540 1152 1552
rect 1174 1540 1181 1552
rect 1117 1392 1124 1404
rect 1145 1392 1152 1404
rect 1174 1392 1181 1404
rect 1117 1191 1124 1203
rect 1145 1191 1152 1203
rect 1174 1191 1181 1203
<< nsubstratencontact >>
rect 1119 1466 1126 1478
rect 1144 1466 1151 1478
rect 1182 1466 1189 1478
rect 1119 1319 1126 1330
rect 1144 1319 1151 1330
rect 1182 1319 1189 1330
rect 1119 1117 1126 1129
rect 1144 1117 1151 1129
rect 1182 1117 1189 1129
use datapathL  datapathL_0
array 0 7 110 0 0 1803
timestamp 1428437267
transform 1 0 30 0 1 562
box 0 -542 110 1261
use rego  rego_2
timestamp 1428352843
transform 1 0 993 0 -1 1840
box 0 -160 110 279
use rego  rego_3
timestamp 1428352843
transform 1 0 1103 0 -1 1840
box 0 -160 110 279
use rego  rego_5
timestamp 1428352843
transform 1 0 1213 0 -1 1840
box 0 -160 110 279
use rego  rego_6
timestamp 1428352843
transform 1 0 1323 0 -1 1840
box 0 -160 110 279
use rego  rego_7
timestamp 1428352843
transform 1 0 1433 0 -1 1840
box 0 -160 110 279
use rego  rego_8
timestamp 1428352843
transform 1 0 1543 0 -1 1840
box 0 -160 110 279
use rego  rego_4
timestamp 1428352843
transform 1 0 993 0 1 1275
box 0 -160 110 279
use rego  rego_1
timestamp 1428352843
transform 1 0 1213 0 1 1275
box 0 -160 110 279
use rego  rego_0
timestamp 1428352843
transform 1 0 1323 0 1 1275
box 0 -160 110 279
use and  and_0
timestamp 1427941063
transform 1 0 1736 0 1 1385
box -25 -23 14 33
use smlogic  smlogic_0
timestamp 1428618667
transform 1 0 1304 0 1 1193
box 123 -146 548 366
use datapathS  datapathS_0
array 0 7 110 0 0 974
timestamp 1428358217
transform 1 0 910 0 1 562
box 0 -542 110 432
<< labels >>
rlabel metal2 1790 495 1815 499 0 INBIT
rlabel metal1 -34 20 4 1822 0 Vdd
rlabel metal1 1828 19 1865 1021 0 GND
rlabel metal1 1140 1423 1157 1437 0 REGMEM
rlabel polysilicon 1203 1229 1208 1249 0 RST
rlabel metal2 1154 1115 1167 1141 0 REGOUT
rlabel metal1 1130 1232 1163 1238 0 REGOUTn
rlabel metal1 1165 1349 1177 1386 0 INCLKn
rlabel metal1 1128 1338 1143 1372 0 INCLK
rlabel polysilicon 1185 1362 1197 1372 0 CLK
rlabel space 1115 1508 1124 1554 0 REGIN
rlabel space 1594 1974 1607 2004 1 valid
rlabel metal1 1696 1423 1704 2014 1 CLK
rlabel metal2 920 1643 928 2006 1 clk
rlabel space 1753 1119 1766 1121 1 start
rlabel metal2 1751 1135 1865 1139 1 start
rlabel space 1844 1028 1852 1344 1 reset
rlabel m2contact 1844 1344 1852 1352 1 reset
rlabel space 1594 1974 1607 2033 1 valid
rlabel space 1594 1974 1607 2029 1 valid
rlabel m2contact 1594 2029 1607 2033 5 valid
rlabel space 813 1785 819 1864 1 divisorin_0
rlabel m2contact 813 1828 819 1833 1 divisorin_0
rlabel m2contact 703 1828 709 1833 1 divisorin_1
rlabel m2contact 593 1828 599 1833 1 divisorin_2
rlabel m2contact 483 1829 489 1834 1 divisorin_3
rlabel m2contact 373 1829 379 1834 1 divisorin_4
rlabel m2contact 263 1828 269 1833 1 divisorin_5
rlabel m2contact 153 1829 159 1834 1 divisorin_6
rlabel metal2 1774 1032 1869 1036 1 dividendin_0
rlabel metal2 1665 1040 1869 1044 1 dividendin_1
rlabel metal2 1555 1048 1869 1052 1 dividendin_2
rlabel metal2 1445 1056 1869 1060 1 dividendin_3
rlabel metal2 1335 1064 1869 1068 1 dividendin_4
rlabel metal2 1225 1072 1869 1076 1 dividendin_5
rlabel metal2 1115 1080 1869 1084 1 dividendin_6
rlabel metal2 1005 1088 1869 1092 1 dividendin_7
rlabel space 1731 -21 1744 46 1 quotient_0
rlabel m2contact 1731 11 1744 17 1 quotient_0
rlabel m2contact 1621 11 1634 17 1 quotient_1
rlabel m2contact 1511 11 1524 17 1 quotient_2
rlabel m2contact 1401 11 1414 17 1 quotient_3
rlabel m2contact 1291 11 1304 17 1 quotient_4
rlabel m2contact 1181 11 1194 17 1 quotient_5
rlabel m2contact 1071 11 1084 17 1 quotient_6
rlabel m2contact 961 11 974 17 1 quotient_7
rlabel m2contact 81 11 94 17 1 remainder_6
rlabel m2contact 191 11 204 17 1 remainder_5
rlabel m2contact 301 11 314 17 1 remainder_4
rlabel m2contact 411 11 424 17 1 remainder_3
rlabel m2contact 521 11 534 17 1 remainder_2
rlabel m2contact 631 11 644 17 1 remainder_1
rlabel m2contact 741 11 754 17 1 remainder_0
rlabel space 1740 1329 1742 1370 1 SB1
rlabel polysilicon 1740 1410 1742 1434 1 SB1
rlabel polysilicon 1730 1410 1732 1434 1 SB0
rlabel polysilicon 1707 1433 1715 1434 1 sign
rlabel space 1613 1113 1651 1115 1 SB0_out
<< end >>
