magic
tech scmos
timestamp 1428611785
<< pwell >>
rect 125 322 139 356
rect 123 177 139 233
rect 452 121 480 150
rect 385 87 480 121
rect 385 71 475 87
rect 123 -24 139 58
rect 385 -26 475 -4
rect 385 -44 480 -26
rect 452 -73 480 -44
<< nwell >>
rect 123 239 139 316
rect 123 64 139 171
rect 385 125 449 155
rect 385 0 475 67
rect 123 -78 139 -30
rect 385 -78 448 -48
<< polysilicon >>
rect 449 149 472 151
rect 449 148 451 149
rect 460 148 462 149
rect 470 148 472 149
rect 406 146 408 148
rect 416 146 418 148
rect 426 146 428 148
rect 436 146 438 148
rect 406 126 408 128
rect 397 121 408 126
rect 416 125 418 128
rect 417 121 418 125
rect 406 118 408 121
rect 416 118 418 121
rect 426 118 428 128
rect 436 118 438 128
rect 406 96 408 98
rect 416 96 418 98
rect 406 84 408 86
rect 416 84 418 86
rect 426 84 428 98
rect 436 84 438 98
rect 460 96 462 108
rect 470 96 472 108
rect 445 86 456 88
rect 406 64 408 74
rect 416 72 418 74
rect 426 72 428 74
rect 416 70 428 72
rect 416 64 418 70
rect 426 64 428 70
rect 436 64 438 74
rect 445 67 447 86
rect 454 84 456 86
rect 464 84 466 86
rect 454 64 456 74
rect 464 64 466 74
rect 406 38 408 44
rect 416 42 418 44
rect 398 36 408 38
rect 398 30 400 36
rect 426 30 428 44
rect 398 26 399 30
rect 427 26 428 30
rect 398 23 400 26
rect 416 23 418 25
rect 426 23 428 26
rect 436 30 438 44
rect 454 42 456 44
rect 464 30 466 44
rect 436 26 437 30
rect 465 26 466 30
rect 436 23 438 26
rect 446 23 448 25
rect 464 23 466 26
rect 398 -7 400 3
rect 416 0 418 3
rect 407 -4 418 0
rect 416 -7 418 -4
rect 426 -7 428 3
rect 436 -7 438 3
rect 446 0 448 3
rect 446 -4 457 0
rect 446 -7 448 -4
rect 464 -7 466 3
rect 398 -19 400 -17
rect 416 -19 418 -17
rect 416 -31 418 -29
rect 426 -31 428 -17
rect 436 -31 438 -17
rect 446 -19 448 -17
rect 464 -19 466 -17
rect 460 -31 462 -29
rect 470 -31 472 -29
rect 416 -44 418 -41
rect 417 -48 418 -44
rect 416 -51 418 -48
rect 426 -51 428 -41
rect 436 -51 438 -41
rect 416 -78 418 -69
rect 426 -81 428 -69
rect 436 -88 438 -69
rect 449 -72 451 -71
rect 460 -72 462 -71
rect 470 -72 472 -71
rect 449 -74 472 -72
rect 429 -91 438 -88
<< ndiffusion >>
rect 404 98 406 118
rect 408 98 410 118
rect 414 98 416 118
rect 418 98 426 118
rect 428 98 436 118
rect 438 98 440 118
rect 458 108 460 148
rect 462 108 464 148
rect 468 108 470 148
rect 472 108 474 148
rect 404 74 406 84
rect 408 74 416 84
rect 418 74 420 84
rect 424 74 426 84
rect 428 74 430 84
rect 434 74 436 84
rect 438 74 440 84
rect 452 74 454 84
rect 456 74 458 84
rect 462 74 464 84
rect 466 74 468 84
rect 396 -17 398 -7
rect 400 -17 402 -7
rect 414 -17 416 -7
rect 418 -17 420 -7
rect 424 -17 426 -7
rect 428 -17 430 -7
rect 434 -17 436 -7
rect 438 -17 440 -7
rect 444 -17 446 -7
rect 448 -17 450 -7
rect 462 -17 464 -7
rect 466 -17 468 -7
rect 414 -41 416 -31
rect 418 -41 426 -31
rect 428 -41 436 -31
rect 438 -41 440 -31
rect 458 -71 460 -31
rect 462 -71 464 -31
rect 468 -71 470 -31
rect 472 -71 474 -31
<< pdiffusion >>
rect 404 128 406 146
rect 408 128 410 146
rect 414 128 416 146
rect 418 128 420 146
rect 424 128 426 146
rect 428 128 430 146
rect 434 128 436 146
rect 438 128 440 146
rect 404 44 406 64
rect 408 44 410 64
rect 414 44 416 64
rect 418 44 420 64
rect 424 44 426 64
rect 428 44 436 64
rect 438 44 440 64
rect 452 44 454 64
rect 456 44 458 64
rect 462 44 464 64
rect 466 44 468 64
rect 396 3 398 23
rect 400 3 402 23
rect 414 3 416 23
rect 418 3 420 23
rect 424 3 426 23
rect 428 3 430 23
rect 434 3 436 23
rect 438 3 440 23
rect 444 3 446 23
rect 448 3 450 23
rect 462 3 464 23
rect 466 3 468 23
rect 414 -69 416 -51
rect 418 -69 420 -51
rect 424 -69 426 -51
rect 428 -69 430 -51
rect 434 -69 436 -51
rect 438 -69 440 -51
<< metal1 >>
rect 128 360 135 362
rect 84 346 135 360
rect 84 213 98 346
rect 128 345 135 346
rect 128 286 134 287
rect 117 272 134 286
rect 128 271 134 272
rect 84 199 134 213
rect 84 12 98 199
rect 128 197 134 199
rect 347 173 376 179
rect 347 169 488 173
rect 368 165 488 169
rect 484 163 488 165
rect 362 161 424 162
rect 358 158 424 161
rect 358 157 365 158
rect 354 145 358 149
rect 378 151 386 155
rect 378 145 382 151
rect 396 151 413 155
rect 410 146 414 151
rect 354 142 360 145
rect 104 138 137 139
rect 104 123 105 138
rect 117 123 137 138
rect 356 122 360 142
rect 369 141 382 145
rect 379 128 393 132
rect 420 146 424 158
rect 484 155 532 163
rect 434 151 475 155
rect 430 146 434 151
rect 447 143 451 144
rect 444 128 454 133
rect 379 122 383 128
rect 400 125 404 128
rect 420 125 424 128
rect 440 125 454 128
rect 356 118 383 122
rect 393 120 397 121
rect 400 121 413 125
rect 420 124 454 125
rect 420 121 449 124
rect 400 118 404 121
rect 440 118 449 121
rect 349 102 373 110
rect 349 33 357 102
rect 444 117 449 118
rect 453 117 454 124
rect 444 108 454 117
rect 478 117 479 126
rect 410 95 414 98
rect 464 95 468 108
rect 381 94 475 95
rect 381 88 397 94
rect 420 88 457 94
rect 471 88 475 94
rect 381 87 475 88
rect 420 84 424 87
rect 440 84 444 87
rect 458 84 462 87
rect 400 71 404 74
rect 430 71 434 74
rect 448 71 452 74
rect 400 67 410 71
rect 434 67 441 71
rect 410 64 414 67
rect 440 64 444 67
rect 448 64 452 67
rect 468 71 472 74
rect 468 67 475 71
rect 468 64 472 67
rect 400 41 404 44
rect 420 41 424 44
rect 458 41 462 44
rect 369 40 475 41
rect 369 33 442 40
rect 463 33 475 40
rect 129 25 134 33
rect 348 25 357 33
rect 392 23 396 33
rect 403 26 409 30
rect 422 26 423 30
rect 430 23 434 33
rect 441 26 442 30
rect 460 26 461 30
rect 468 23 472 33
rect 84 -2 145 12
rect 84 -5 98 -2
rect 128 -4 134 -2
rect 348 -4 373 12
rect 406 3 407 23
rect 403 0 407 3
rect 410 0 414 3
rect 450 0 454 3
rect 410 -4 420 0
rect 403 -7 407 -4
rect 420 -7 424 -4
rect 444 -4 454 0
rect 457 3 458 23
rect 457 0 461 3
rect 472 -4 475 0
rect 440 -7 444 -4
rect 457 -7 461 -4
rect 406 -17 407 -7
rect 457 -17 458 -7
rect 392 -20 396 -17
rect 410 -20 414 -17
rect 430 -20 434 -17
rect 450 -20 454 -17
rect 468 -20 472 -17
rect 381 -21 475 -20
rect 381 -27 395 -21
rect 420 -27 475 -21
rect 381 -28 475 -27
rect 410 -31 414 -28
rect 464 -31 468 -28
rect 444 -41 454 -31
rect 440 -44 449 -41
rect 397 -48 413 -44
rect 424 -48 449 -44
rect 453 -48 454 -41
rect 420 -51 424 -48
rect 440 -51 454 -48
rect 128 -63 134 -62
rect 106 -66 139 -63
rect 115 -77 139 -66
rect 106 -79 139 -77
rect 346 -78 361 -62
rect 447 -67 451 -66
rect 410 -74 414 -69
rect 430 -74 434 -69
rect 478 -48 479 -41
rect 369 -78 387 -74
rect 406 -78 475 -74
rect 197 -85 287 -81
rect 307 -85 425 -81
rect 283 -88 287 -85
rect 283 -92 425 -88
rect 524 -115 532 155
rect 540 -146 548 151
<< metal2 >>
rect 148 363 366 366
rect 148 358 154 363
rect 258 352 358 358
rect 105 138 116 272
rect 354 161 358 352
rect 362 153 366 363
rect 383 168 484 169
rect 383 164 485 168
rect 358 149 366 153
rect 373 161 485 164
rect 373 156 383 161
rect 481 159 485 161
rect 373 151 382 156
rect 417 151 430 155
rect 481 151 540 159
rect 363 130 369 141
rect 105 -66 116 123
rect 115 -77 116 -66
rect 361 41 369 130
rect 373 110 381 151
rect 385 139 447 140
rect 385 136 451 139
rect 361 -62 369 33
rect 373 12 381 87
rect 373 -20 381 -4
rect 385 -52 389 136
rect 464 132 480 135
rect 397 128 405 132
rect 393 -44 397 116
rect 401 -39 405 128
rect 410 131 480 132
rect 410 128 468 131
rect 410 71 414 128
rect 453 117 479 124
rect 430 108 481 112
rect 430 71 434 108
rect 448 63 475 67
rect 409 34 446 38
rect 409 30 413 34
rect 442 30 446 34
rect 418 22 422 26
rect 456 22 460 26
rect 418 18 460 22
rect 444 -4 468 0
rect 420 -31 424 -4
rect 420 -35 483 -31
rect 401 -43 424 -39
rect 420 -44 424 -43
rect 453 -48 479 -41
rect 385 -56 451 -52
rect 184 -81 197 -77
rect 294 -81 307 -76
rect 447 -62 451 -56
<< ntransistor >>
rect 406 98 408 118
rect 416 98 418 118
rect 426 98 428 118
rect 436 98 438 118
rect 460 108 462 148
rect 470 108 472 148
rect 406 74 408 84
rect 416 74 418 84
rect 426 74 428 84
rect 436 74 438 84
rect 454 74 456 84
rect 464 74 466 84
rect 398 -17 400 -7
rect 416 -17 418 -7
rect 426 -17 428 -7
rect 436 -17 438 -7
rect 446 -17 448 -7
rect 464 -17 466 -7
rect 416 -41 418 -31
rect 426 -41 428 -31
rect 436 -41 438 -31
rect 460 -71 462 -31
rect 470 -71 472 -31
<< ptransistor >>
rect 406 128 408 146
rect 416 128 418 146
rect 426 128 428 146
rect 436 128 438 146
rect 406 44 408 64
rect 416 44 418 64
rect 426 44 428 64
rect 436 44 438 64
rect 454 44 456 64
rect 464 44 466 64
rect 398 3 400 23
rect 416 3 418 23
rect 426 3 428 23
rect 436 3 438 23
rect 446 3 448 23
rect 464 3 466 23
rect 416 -69 418 -51
rect 426 -69 428 -51
rect 436 -69 438 -51
<< polycontact >>
rect 447 144 451 148
rect 393 121 397 125
rect 413 121 417 125
rect 441 67 445 71
rect 399 26 403 30
rect 423 26 427 30
rect 437 26 441 30
rect 461 26 465 30
rect 403 -4 407 0
rect 457 -4 461 0
rect 413 -48 417 -44
rect 425 -85 429 -81
rect 447 -71 451 -67
rect 425 -92 429 -88
<< ndcontact >>
rect 400 98 404 118
rect 410 98 414 118
rect 440 98 444 118
rect 454 108 458 148
rect 464 108 468 148
rect 474 108 478 148
rect 400 74 404 84
rect 420 74 424 84
rect 430 74 434 84
rect 440 74 444 84
rect 448 74 452 84
rect 458 74 462 84
rect 468 74 472 84
rect 392 -17 396 -7
rect 402 -17 406 -7
rect 410 -17 414 -7
rect 420 -17 424 -7
rect 430 -17 434 -7
rect 440 -17 444 -7
rect 450 -17 454 -7
rect 458 -17 462 -7
rect 468 -17 472 -7
rect 410 -41 414 -31
rect 440 -41 444 -31
rect 454 -71 458 -31
rect 464 -71 468 -31
rect 474 -71 478 -31
<< pdcontact >>
rect 400 128 404 146
rect 410 128 414 146
rect 420 128 424 146
rect 430 128 434 146
rect 440 128 444 146
rect 400 44 404 64
rect 410 44 414 64
rect 420 44 424 64
rect 440 44 444 64
rect 448 44 452 64
rect 458 44 462 64
rect 468 44 472 64
rect 392 3 396 23
rect 402 3 406 23
rect 410 3 414 23
rect 420 3 424 23
rect 430 3 434 23
rect 440 3 444 23
rect 450 3 454 23
rect 458 3 462 23
rect 468 3 472 23
rect 410 -69 414 -51
rect 420 -69 424 -51
rect 430 -69 434 -51
rect 440 -69 444 -51
<< m2contact >>
rect 105 272 117 287
rect 354 157 358 161
rect 354 149 358 153
rect 413 151 417 155
rect 105 123 117 138
rect 363 141 369 145
rect 393 128 397 132
rect 430 151 434 155
rect 447 139 451 143
rect 393 116 397 120
rect 373 102 381 110
rect 449 117 453 124
rect 479 117 483 126
rect 373 87 381 95
rect 410 67 414 71
rect 430 67 434 71
rect 448 67 452 71
rect 361 33 369 41
rect 409 26 413 30
rect 418 26 422 30
rect 442 26 446 30
rect 456 26 460 30
rect 373 -4 381 12
rect 420 -4 424 0
rect 440 -4 444 0
rect 468 -4 472 0
rect 373 -28 381 -20
rect 393 -48 397 -44
rect 420 -48 424 -44
rect 449 -48 453 -41
rect 105 -77 115 -66
rect 361 -78 369 -62
rect 447 -66 451 -62
rect 479 -48 483 -41
rect 184 -85 197 -81
rect 294 -85 307 -81
rect 540 151 548 159
<< psubstratepcontact >>
rect 397 88 420 94
rect 457 88 471 94
rect 395 -27 420 -21
<< nsubstratencontact >>
rect 386 148 396 155
rect 442 33 463 40
rect 387 -78 406 -74
use rego  rego_0
timestamp 1428352843
transform 1 0 133 0 1 82
box 0 -160 110 279
use rego  rego_1
timestamp 1428352843
transform 1 0 243 0 1 82
box 0 -160 110 279
<< labels >>
rlabel metal2 385 -56 451 -52 1 start
rlabel metal1 420 -48 444 -44 1 nextSB1
rlabel metal2 374 -28 380 95 3 Gnd
rlabel polysilicon 436 -81 438 -71 1 SB1
rlabel polysilicon 426 -81 428 -71 1 SB0
rlabel metal1 397 -48 413 -44 1 sign
rlabel metal1 472 -4 475 0 7 add
rlabel metal2 448 63 475 67 1 sel0
rlabel metal1 468 64 472 74 1 sel1
rlabel metal2 401 -43 424 -39 1 nextSB1
rlabel metal1 347 169 376 179 1 clk
rlabel metal1 540 -146 548 151 7 reset
rlabel metal2 420 -35 483 -31 1 inbit
rlabel metal2 361 41 369 141 3 Vdd
rlabel metal2 430 108 481 112 1 load
rlabel metal2 464 131 480 135 1 shift
rlabel metal1 420 146 424 162 1 nextSB0
rlabel metal1 420 121 444 125 1 nextSB0
<< end >>
